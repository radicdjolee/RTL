----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/10/2022 10:08:27 PM
-- Design Name: 
-- Module Name: cos_rom - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cos_rom is
    generic (
	       WIDTH : integer := 32;
	       WIDTH_2 : integer := 64;
	       WIDTH_3 : integer := 96; 
	       WADDR   : integer := 10
    );
    port(
        address_cos_0 : in  std_logic_vector(WADDR-1 downto 0);
        dout_cos_0    : out std_logic_vector(WIDTH-1 downto 0)
    );
end cos_rom;

architecture Behavioral of cos_rom is
  type mem is array ( 0 to 647) of std_logic_vector(WIDTH-1 downto 0);
  constant my_Rom : mem := (

0 => "00111111001011001111001101110111",
1 => "10111111010010110001100100101111",
2 => "10111111000010011000110001111110",
3 => "00111111011000110001001100100111",
4 => "00111110110000111110111100000111",
5 => "10111111011101000010011011001100",
6 => "10111110010111011010001001110011",
7 => "00111111011111011100111101010111",
8 => "00111101001100101010101001000010",
9 => "10111111011111111100000110011100",
10 => "00111110000001011010100010011100",
11 => "00111111011110011110111010001001",
12 => "10111110100110011111011000100011",
13 => "10111111011011001000001101100110",
14 => "00111110111011000110101001011101",
15 => "00111111010101111110100001111001",
16 => "10111111000110111101011111000011",
17 => "10111111001111001011111000101111",
18 => "00111111000110111101011111000011",
19 => "10111111011011001000001101100110",
20 => "10111110000001011010100010011100",
21 => "00111111011111011100111101010111",
22 => "10111110110000111110111100000111",
23 => "10111111010010110001100100101111",
24 => "00111111010010110001100100101111",
25 => "00111110110000111110111100000111",
26 => "10111111011111011100111101010111",
27 => "00111110000001011010100010011100",
28 => "00111111011011001000001101100110",
29 => "10111111000110111101011111000011",
30 => "10111111000110111101011111000011",
31 => "00111111011011001000001101100110",
32 => "00111110000001011010100010011100",
33 => "10111111011111011100111101010111",
34 => "00111110110000111110111100000111",
35 => "00111111010010110001100100101111",
36 => "00111111000010011000110001111110",
37 => "10111111011111011100111101010111",
38 => "00111110100110011111011000100011",
39 => "00111111001111001011111000101111",
40 => "10111111011011001000001101100110",
41 => "00111101001100101010101001000010",
42 => "00111111011000110001001100100111",
43 => "10111111010010110001100100101111",
44 => "10111110010111011010001001110011",
45 => "00111111011110011110111010001001",
46 => "10111111000110111101011111000011",
47 => "10111110111011000110101001011101",
48 => "00111111011111111100000110011100",
49 => "10111110110000111110111100000111",
50 => "10111111001011001111001101110111",
51 => "00111111011101000010011011001100",
52 => "10111110000001011010100010011100",
53 => "10111111010101111110100001111001",
54 => "00111110111011000110101001011101",
55 => "10111111011111011100111101010111",
56 => "00111111001011001111001101110111",
57 => "00111110010111011010001001110011",
58 => "10111111011011001000001101100110",
59 => "00111111010101111110100001111001",
60 => "10111101001100101010101001000010",
61 => "10111111010010110001100100101111",
62 => "00111111011101000010011011001100",
63 => "10111110100110011111011000100011",
64 => "10111111000110111101011111000011",
65 => "00111111011111111100000110011100",
66 => "10111111000010011000110001111110",
67 => "10111110110000111110111100000111",
68 => "00111111011110011110111010001001",
69 => "10111111001111001011111000101111",
70 => "10111110000001011010100010011100",
71 => "00111111011000110001001100100111",
72 => "00111110110000111110111100000111",
73 => "10111111011011001000001101100110",
74 => "00111111011011001000001101100110",
75 => "10111110110000111110111100000111",
76 => "10111110110000111110111100000111",
77 => "00111111011011001000001101100110",
78 => "10111111011011001000001101100110",
79 => "00111110110000111110111100000111",
80 => "00111110110000111110111100000111",
81 => "10111111011011001000001101100110",
82 => "00111111011011001000001101100110",
83 => "10111110110000111110111100000111",
84 => "10111110110000111110111100000111",
85 => "00111111011011001000001101100110",
86 => "10111111011011001000001101100110",
87 => "00111110110000111110111100000111",
88 => "00111110110000111110111100000111",
89 => "10111111011011001000001101100110",
90 => "00111110100110011111011000100011",
91 => "10111111010010110001100100101111",
92 => "00111111011111111100000110011100",
93 => "10111111010101111110100001111001",
94 => "00111110110000111110111100000111",
95 => "00111110010111011010001001110011",
96 => "10111111001111001011111000101111",
97 => "00111111011111011100111101010111",
98 => "10111111011000110001001100100111",
99 => "00111110111011000110101001011101",
100 => "00111110000001011010100010011100",
101 => "10111111001011001111001101110111",
102 => "00111111011110011110111010001001",
103 => "10111111011011001000001101100110",
104 => "00111111000010011000110001111110",
105 => "00111101001100101010101001000010",
106 => "10111111000110111101011111000011",
107 => "00111111011101000010011011001100",
108 => "00111110010111011010001001110011",
109 => "10111111000110111101011111000011",
110 => "00111111011000110001001100100111",
111 => "10111111011111111100000110011100",
112 => "00111111011011001000001101100110",
113 => "10111111001011001111001101110111",
114 => "00111110100110011111011000100011",
115 => "00111110000001011010100010011100",
116 => "10111111000010011000110001111110",
117 => "00111111010101111110100001111001",
118 => "10111111011111011100111101010111",
119 => "00111111011101000010011011001100",
120 => "10111111001111001011111000101111",
121 => "00111110110000111110111100000111",
122 => "00111101001100101010101001000010",
123 => "10111110111011000110101001011101",
124 => "00111111010010110001100100101111",
125 => "10111111011110011110111010001001",
126 => "00111110000001011010100010011100",
127 => "10111110110000111110111100000111",
128 => "00111111000110111101011111000011",
129 => "10111111010010110001100100101111",
130 => "00111111011011001000001101100110",
131 => "10111111011111011100111101010111",
132 => "00111111011111011100111101010111",
133 => "10111111011011001000001101100110",
134 => "00111111010010110001100100101111",
135 => "10111111000110111101011111000011",
136 => "00111110110000111110111100000111",
137 => "10111110000001011010100010011100",
138 => "10111110000001011010100010011100",
139 => "00111110110000111110111100000111",
140 => "10111111000110111101011111000011",
141 => "00111111010010110001100100101111",
142 => "10111111011011001000001101100110",
143 => "00111111011111011100111101010111",
144 => "00111101001100101010101001000010",
145 => "10111110000001011010100010011100",
146 => "00111110010111011010001001110011",
147 => "10111110100110011111011000100011",
148 => "00111110110000111110111100000111",
149 => "10111110111011000110101001011101",
150 => "00111111000010011000110001111110",
151 => "10111111000110111101011111000011",
152 => "00111111001011001111001101110111",
153 => "10111111001111001011111000101111",
154 => "00111111010010110001100100101111",
155 => "10111111010101111110100001111001",
156 => "00111111011000110001001100100111",
157 => "10111111011011001000001101100110",
158 => "00111111011101000010011011001100",
159 => "10111111011110011110111010001001",
160 => "00111111011111011100111101010111",
161 => "10111111011111111100000110011100",
162 => "10111101001100101010101001000010",
163 => "00111110000001011010100010011100",
164 => "10111110010111011010001001110011",
165 => "00111110100110011111011000100011",
166 => "10111110110000111110111100000111",
167 => "00111110111011000110101001011101",
168 => "10111111000010011000110001111110",
169 => "00111111000110111101011111000011",
170 => "10111111001011001111001101110111",
171 => "00111111001111001011111000101111",
172 => "10111111010010110001100100101111",
173 => "00111111010101111110100001111001",
174 => "10111111011000110001001100100111",
175 => "00111111011011001000001101100110",
176 => "10111111011101000010011011001100",
177 => "00111111011110011110111010001001",
178 => "10111111011111011100111101010111",
179 => "00111111011111111100000110011100",
180 => "10111110000001011010100010011100",
181 => "00111110110000111110111100000111",
182 => "10111111000110111101011111000011",
183 => "00111111010010110001100100101111",
184 => "10111111011011001000001101100110",
185 => "00111111011111011100111101010111",
186 => "10111111011111011100111101010111",
187 => "00111111011011001000001101100110",
188 => "10111111010010110001100100101111",
189 => "00111111000110111101011111000011",
190 => "10111110110000111110111100000111",
191 => "00111110000001011010100010011100",
192 => "00111110000001011010100010011100",
193 => "10111110110000111110111100000111",
194 => "00111111000110111101011111000011",
195 => "10111111010010110001100100101111",
196 => "00111111011011001000001101100110",
197 => "10111111011111011100111101010111",
198 => "10111110010111011010001001110011",
199 => "00111111000110111101011111000011",
200 => "10111111011000110001001100100111",
201 => "00111111011111111100000110011100",
202 => "10111111011011001000001101100110",
203 => "00111111001011001111001101110111",
204 => "10111110100110011111011000100011",
205 => "10111110000001011010100010011100",
206 => "00111111000010011000110001111110",
207 => "10111111010101111110100001111001",
208 => "00111111011111011100111101010111",
209 => "10111111011101000010011011001100",
210 => "00111111001111001011111000101111",
211 => "10111110110000111110111100000111",
212 => "10111101001100101010101001000010",
213 => "00111110111011000110101001011101",
214 => "10111111010010110001100100101111",
215 => "00111111011110011110111010001001",
216 => "10111110100110011111011000100011",
217 => "00111111010010110001100100101111",
218 => "10111111011111111100000110011100",
219 => "00111111010101111110100001111001",
220 => "10111110110000111110111100000111",
221 => "10111110010111011010001001110011",
222 => "00111111001111001011111000101111",
223 => "10111111011111011100111101010111",
224 => "00111111011000110001001100100111",
225 => "10111110111011000110101001011101",
226 => "10111110000001011010100010011100",
227 => "00111111001011001111001101110111",
228 => "10111111011110011110111010001001",
229 => "00111111011011001000001101100110",
230 => "10111111000010011000110001111110",
231 => "10111101001100101010101001000010",
232 => "00111111000110111101011111000011",
233 => "10111111011101000010011011001100",
234 => "10111110110000111110111100000111",
235 => "00111111011011001000001101100110",
236 => "10111111011011001000001101100110",
237 => "00111110110000111110111100000111",
238 => "00111110110000111110111100000111",
239 => "10111111011011001000001101100110",
240 => "00111111011011001000001101100110",
241 => "10111110110000111110111100000111",
242 => "10111110110000111110111100000111",
243 => "00111111011011001000001101100110",
244 => "10111111011011001000001101100110",
245 => "00111110110000111110111100000111",
246 => "00111110110000111110111100000111",
247 => "10111111011011001000001101100110",
248 => "00111111011011001000001101100110",
249 => "10111110110000111110111100000111",
250 => "10111110110000111110111100000111",
251 => "00111111011011001000001101100110",
252 => "10111110111011000110101001011101",
253 => "00111111011111011100111101010111",
254 => "10111111001011001111001101110111",
255 => "10111110010111011010001001110011",
256 => "00111111011011001000001101100110",
257 => "10111111010101111110100001111001",
258 => "00111101001100101010101001000010",
259 => "00111111010010110001100100101111",
260 => "10111111011101000010011011001100",
261 => "00111110100110011111011000100011",
262 => "00111111000110111101011111000011",
263 => "10111111011111111100000110011100",
264 => "00111111000010011000110001111110",
265 => "00111110110000111110111100000111",
266 => "10111111011110011110111010001001",
267 => "00111111001111001011111000101111",
268 => "00111110000001011010100010011100",
269 => "10111111011000110001001100100111",
270 => "10111111000010011000110001111110",
271 => "00111111011111011100111101010111",
272 => "10111110100110011111011000100011",
273 => "10111111001111001011111000101111",
274 => "00111111011011001000001101100110",
275 => "10111101001100101010101001000010",
276 => "10111111011000110001001100100111",
277 => "00111111010010110001100100101111",
278 => "00111110010111011010001001110011",
279 => "10111111011110011110111010001001",
280 => "00111111000110111101011111000011",
281 => "00111110111011000110101001011101",
282 => "10111111011111111100000110011100",
283 => "00111110110000111110111100000111",
284 => "00111111001011001111001101110111",
285 => "10111111011101000010011011001100",
286 => "00111110000001011010100010011100",
287 => "00111111010101111110100001111001",
288 => "10111111000110111101011111000011",
289 => "00111111011011001000001101100110",
290 => "00111110000001011010100010011100",
291 => "10111111011111011100111101010111",
292 => "00111110110000111110111100000111",
293 => "00111111010010110001100100101111",
294 => "10111111010010110001100100101111",
295 => "10111110110000111110111100000111",
296 => "00111111011111011100111101010111",
297 => "10111110000001011010100010011100",
298 => "10111111011011001000001101100110",
299 => "00111111000110111101011111000011",
300 => "00111111000110111101011111000011",
301 => "10111111011011001000001101100110",
302 => "10111110000001011010100010011100",
303 => "00111111011111011100111101010111",
304 => "10111110110000111110111100000111",
305 => "10111111010010110001100100101111",
306 => "10111111001011001111001101110111",
307 => "00111111010010110001100100101111",
308 => "00111111000010011000110001111110",
309 => "10111111011000110001001100100111",
310 => "10111110110000111110111100000111",
311 => "00111111011101000010011011001100",
312 => "00111110010111011010001001110011",
313 => "10111111011111011100111101010111",
314 => "10111101001100101010101001000010",
315 => "00111111011111111100000110011100",
316 => "10111110000001011010100010011100",
317 => "10111111011110011110111010001001",
318 => "00111110100110011111011000100011",
319 => "00111111011011001000001101100110",
320 => "10111110111011000110101001011101",
321 => "10111111010101111110100001111001",
322 => "00111111000110111101011111000011",
323 => "00111111001111001011111000101111",
324 => "10111111001111001011111000101111",
325 => "00111111000110111101011111000011",
326 => "00111111010101111110100001111001",
327 => "10111110111011000110101001011101",
328 => "10111111011011001000001101100110",
329 => "00111110100110011111011000100011",
330 => "00111111011110011110111010001001",
331 => "10111110000001011010100010011100",
332 => "10111111011111111100000110011100",
333 => "10111101001100101010101001000010",
334 => "00111111011111011100111101010111",
335 => "00111110010111011010001001110011",
336 => "10111111011101000010011011001100",
337 => "10111110110000111110111100000111",
338 => "00111111011000110001001100100111",
339 => "00111111000010011000110001111110",
340 => "10111111010010110001100100101111",
341 => "10111111001011001111001101110111",
342 => "10111111010010110001100100101111",
343 => "00111110110000111110111100000111",
344 => "00111111011111011100111101010111",
345 => "00111110000001011010100010011100",
346 => "10111111011011001000001101100110",
347 => "10111111000110111101011111000011",
348 => "00111111000110111101011111000011",
349 => "00111111011011001000001101100110",
350 => "10111110000001011010100010011100",
351 => "10111111011111011100111101010111",
352 => "10111110110000111110111100000111",
353 => "00111111010010110001100100101111",
354 => "00111111010010110001100100101111",
355 => "10111110110000111110111100000111",
356 => "10111111011111011100111101010111",
357 => "10111110000001011010100010011100",
358 => "00111111011011001000001101100110",
359 => "00111111000110111101011111000011",
360 => "10111111010101111110100001111001",
361 => "00111110000001011010100010011100",
362 => "00111111011101000010011011001100",
363 => "00111111001011001111001101110111",
364 => "10111110110000111110111100000111",
365 => "10111111011111111100000110011100",
366 => "10111110111011000110101001011101",
367 => "00111111000110111101011111000011",
368 => "00111111011110011110111010001001",
369 => "00111110010111011010001001110011",
370 => "10111111010010110001100100101111",
371 => "10111111011000110001001100100111",
372 => "00111101001100101010101001000010",
373 => "00111111011011001000001101100110",
374 => "00111111001111001011111000101111",
375 => "10111110100110011111011000100011",
376 => "10111111011111011100111101010111",
377 => "10111111000010011000110001111110",
378 => "10111111011000110001001100100111",
379 => "10111110000001011010100010011100",
380 => "00111111001111001011111000101111",
381 => "00111111011110011110111010001001",
382 => "00111110110000111110111100000111",
383 => "10111111000010011000110001111110",
384 => "10111111011111111100000110011100",
385 => "10111111000110111101011111000011",
386 => "00111110100110011111011000100011",
387 => "00111111011101000010011011001100",
388 => "00111111010010110001100100101111",
389 => "10111101001100101010101001000010",
390 => "10111111010101111110100001111001",
391 => "10111111011011001000001101100110",
392 => "10111110010111011010001001110011",
393 => "00111111001011001111001101110111",
394 => "00111111011111011100111101010111",
395 => "00111110111011000110101001011101",
396 => "10111111011011001000001101100110",
397 => "10111110110000111110111100000111",
398 => "00111110110000111110111100000111",
399 => "00111111011011001000001101100110",
400 => "00111111011011001000001101100110",
401 => "00111110110000111110111100000111",
402 => "10111110110000111110111100000111",
403 => "10111111011011001000001101100110",
404 => "10111111011011001000001101100110",
405 => "10111110110000111110111100000111",
406 => "00111110110000111110111100000111",
407 => "00111111011011001000001101100110",
408 => "00111111011011001000001101100110",
409 => "00111110110000111110111100000111",
410 => "10111110110000111110111100000111",
411 => "10111111011011001000001101100110",
412 => "10111111011011001000001101100110",
413 => "10111110110000111110111100000111",
414 => "10111111011101000010011011001100",
415 => "10111111000110111101011111000011",
416 => "10111101001100101010101001000010",
417 => "00111111000010011000110001111110",
418 => "00111111011011001000001101100110",
419 => "00111111011110011110111010001001",
420 => "00111111001011001111001101110111",
421 => "00111110000001011010100010011100",
422 => "10111110111011000110101001011101",
423 => "10111111011000110001001100100111",
424 => "10111111011111011100111101010111",
425 => "10111111001111001011111000101111",
426 => "10111110010111011010001001110011",
427 => "00111110110000111110111100000111",
428 => "00111111010101111110100001111001",
429 => "00111111011111111100000110011100",
430 => "00111111010010110001100100101111",
431 => "00111110100110011111011000100011",
432 => "10111111011110011110111010001001",
433 => "10111111010010110001100100101111",
434 => "10111110111011000110101001011101",
435 => "10111101001100101010101001000010",
436 => "00111110110000111110111100000111",
437 => "00111111001111001011111000101111",
438 => "00111111011101000010011011001100",
439 => "00111111011111011100111101010111",
440 => "00111111010101111110100001111001",
441 => "00111111000010011000110001111110",
442 => "00111110000001011010100010011100",
443 => "10111110100110011111011000100011",
444 => "10111111001011001111001101110111",
445 => "10111111011011001000001101100110",
446 => "10111111011111111100000110011100",
447 => "10111111011000110001001100100111",
448 => "10111111000110111101011111000011",
449 => "10111110010111011010001001110011",
450 => "10111111011111011100111101010111",
451 => "10111111011011001000001101100110",
452 => "10111111010010110001100100101111",
453 => "10111111000110111101011111000011",
454 => "10111110110000111110111100000111",
455 => "10111110000001011010100010011100",
456 => "00111110000001011010100010011100",
457 => "00111110110000111110111100000111",
458 => "00111111000110111101011111000011",
459 => "00111111010010110001100100101111",
460 => "00111111011011001000001101100110",
461 => "00111111011111011100111101010111",
462 => "00111111011111011100111101010111",
463 => "00111111011011001000001101100110",
464 => "00111111010010110001100100101111",
465 => "00111111000110111101011111000011",
466 => "00111110110000111110111100000111",
467 => "00111110000001011010100010011100",
468 => "10111111011111111100000110011100",
469 => "10111111011111011100111101010111",
470 => "10111111011110011110111010001001",
471 => "10111111011101000010011011001100",
472 => "10111111011011001000001101100110",
473 => "10111111011000110001001100100111",
474 => "10111111010101111110100001111001",
475 => "10111111010010110001100100101111",
476 => "10111111001111001011111000101111",
477 => "10111111001011001111001101110111",
478 => "10111111000110111101011111000011",
479 => "10111111000010011000110001111110",
480 => "10111110111011000110101001011101",
481 => "10111110110000111110111100000111",
482 => "10111110100110011111011000100011",
483 => "10111110010111011010001001110011",
484 => "10111110000001011010100010011100",
485 => "10111101001100101010101001000010",
486 => "10111111011111111100000110011100",
487 => "10111111011111011100111101010111",
488 => "10111111011110011110111010001001",
489 => "10111111011101000010011011001100",
490 => "10111111011011001000001101100110",
491 => "10111111011000110001001100100111",
492 => "10111111010101111110100001111001",
493 => "10111111010010110001100100101111",
494 => "10111111001111001011111000101111",
495 => "10111111001011001111001101110111",
496 => "10111111000110111101011111000011",
497 => "10111111000010011000110001111110",
498 => "10111110111011000110101001011101",
499 => "10111110110000111110111100000111",
500 => "10111110100110011111011000100011",
501 => "10111110010111011010001001110011",
502 => "10111110000001011010100010011100",
503 => "10111101001100101010101001000010",
504 => "10111111011111011100111101010111",
505 => "10111111011011001000001101100110",
506 => "10111111010010110001100100101111",
507 => "10111111000110111101011111000011",
508 => "10111110110000111110111100000111",
509 => "10111110000001011010100010011100",
510 => "00111110000001011010100010011100",
511 => "00111110110000111110111100000111",
512 => "00111111000110111101011111000011",
513 => "00111111010010110001100100101111",
514 => "00111111011011001000001101100110",
515 => "00111111011111011100111101010111",
516 => "00111111011111011100111101010111",
517 => "00111111011011001000001101100110",
518 => "00111111010010110001100100101111",
519 => "00111111000110111101011111000011",
520 => "00111110110000111110111100000111",
521 => "00111110000001011010100010011100",
522 => "10111111011110011110111010001001",
523 => "10111111010010110001100100101111",
524 => "10111110111011000110101001011101",
525 => "10111101001100101010101001000010",
526 => "00111110110000111110111100000111",
527 => "00111111001111001011111000101111",
528 => "00111111011101000010011011001100",
529 => "00111111011111011100111101010111",
530 => "00111111010101111110100001111001",
531 => "00111111000010011000110001111110",
532 => "00111110000001011010100010011100",
533 => "10111110100110011111011000100011",
534 => "10111111001011001111001101110111",
535 => "10111111011011001000001101100110",
536 => "10111111011111111100000110011100",
537 => "10111111011000110001001100100111",
538 => "10111111000110111101011111000011",
539 => "10111110010111011010001001110011",
540 => "10111111011101000010011011001100",
541 => "10111111000110111101011111000011",
542 => "10111101001100101010101001000010",
543 => "00111111000010011000110001111110",
544 => "00111111011011001000001101100110",
545 => "00111111011110011110111010001001",
546 => "00111111001011001111001101110111",
547 => "00111110000001011010100010011100",
548 => "10111110111011000110101001011101",
549 => "10111111011000110001001100100111",
550 => "10111111011111011100111101010111",
551 => "10111111001111001011111000101111",
552 => "10111110010111011010001001110011",
553 => "00111110110000111110111100000111",
554 => "00111111010101111110100001111001",
555 => "00111111011111111100000110011100",
556 => "00111111010010110001100100101111",
557 => "00111110100110011111011000100011",
558 => "10111111011011001000001101100110",
559 => "10111110110000111110111100000111",
560 => "00111110110000111110111100000111",
561 => "00111111011011001000001101100110",
562 => "00111111011011001000001101100110",
563 => "00111110110000111110111100000111",
564 => "10111110110000111110111100000111",
565 => "10111111011011001000001101100110",
566 => "10111111011011001000001101100110",
567 => "10111110110000111110111100000111",
568 => "00111110110000111110111100000111",
569 => "00111111011011001000001101100110",
570 => "00111111011011001000001101100110",
571 => "00111110110000111110111100000111",
572 => "10111110110000111110111100000111",
573 => "10111111011011001000001101100110",
574 => "10111111011011001000001101100110",
575 => "10111110110000111110111100000111",
576 => "10111111011000110001001100100111",
577 => "10111110000001011010100010011100",
578 => "00111111001111001011111000101111",
579 => "00111111011110011110111010001001",
580 => "00111110110000111110111100000111",
581 => "10111111000010011000110001111110",
582 => "10111111011111111100000110011100",
583 => "10111111000110111101011111000011",
584 => "00111110100110011111011000100011",
585 => "00111111011101000010011011001100",
586 => "00111111010010110001100100101111",
587 => "10111101001100101010101001000010",
588 => "10111111010101111110100001111001",
589 => "10111111011011001000001101100110",
590 => "10111110010111011010001001110011",
591 => "00111111001011001111001101110111",
592 => "00111111011111011100111101010111",
593 => "00111110111011000110101001011101",
594 => "10111111010101111110100001111001",
595 => "00111110000001011010100010011100",
596 => "00111111011101000010011011001100",
597 => "00111111001011001111001101110111",
598 => "10111110110000111110111100000111",
599 => "10111111011111111100000110011100",
600 => "10111110111011000110101001011101",
601 => "00111111000110111101011111000011",
602 => "00111111011110011110111010001001",
603 => "00111110010111011010001001110011",
604 => "10111111010010110001100100101111",
605 => "10111111011000110001001100100111",
606 => "00111101001100101010101001000010",
607 => "00111111011011001000001101100110",
608 => "00111111001111001011111000101111",
609 => "10111110100110011111011000100011",
610 => "10111111011111011100111101010111",
611 => "10111111000010011000110001111110",
612 => "10111111010010110001100100101111",
613 => "00111110110000111110111100000111",
614 => "00111111011111011100111101010111",
615 => "00111110000001011010100010011100",
616 => "10111111011011001000001101100110",
617 => "10111111000110111101011111000011",
618 => "00111111000110111101011111000011",
619 => "00111111011011001000001101100110",
620 => "10111110000001011010100010011100",
621 => "10111111011111011100111101010111",
622 => "10111110110000111110111100000111",
623 => "00111111010010110001100100101111",
624 => "00111111010010110001100100101111",
625 => "10111110110000111110111100000111",
626 => "10111111011111011100111101010111",
627 => "10111110000001011010100010011100",
628 => "00111111011011001000001101100110",
629 => "00111111000110111101011111000011",
630 => "10111111001111001011111000101111",
631 => "00111111000110111101011111000011",
632 => "00111111010101111110100001111001",
633 => "10111110111011000110101001011101",
634 => "10111111011011001000001101100110",
635 => "00111110100110011111011000100011",
636 => "00111111011110011110111010001001",
637 => "10111110000001011010100010011100",
638 => "10111111011111111100000110011100",
639 => "10111101001100101010101001000010",
640 => "00111111011111011100111101010111",
641 => "00111110010111011010001001110011",
642 => "10111111011101000010011011001100",
643 => "10111110110000111110111100000111",
644 => "00111111011000110001001100100111",
645 => "00111111000010011000110001111110",
646 => "10111111010010110001100100101111",
647 => "10111111001011001111001101110111");
begin

    main : process(address_cos_0)
    begin
        dout_cos_0 <= my_Rom(to_integer(unsigned(address_cos_0)));
    end process main;

end Behavioral;

